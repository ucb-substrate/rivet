module decoder(
  input [3:0] A,
  output [15:0] Z,
  input clk
);

	
// Only one output should ever be high.  For example,
// Z[2] = !A[3] & !A[2] & A[1] & !A[0], etc

// Hint: a 2 to 1 mux looks like:
// assign y = (sel) ? b : a;
// And you can replace "a" with a further condition
// assign y = (sel1) ? c
//          : (sel2) ? b
//          : a
// and sel1 can be a condition like:
// A == 4'd0

assign Z
  = (A[3:0] == 4'b0000) ? 16'b0000_0000_0000_0001
  : (A[3:0] == 4'b0001) ? 16'b0000_0000_0000_0010
  : (A[3:0] == 4'b0010) ? 16'b0000_0000_0000_0100
  : (A[3:0] == 4'b0011) ? 16'b0000_0000_0000_1000
  : (A[3:0] == 4'b0100) ? 16'b0000_0000_0001_0000
  : (A[3:0] == 4'b0101) ? 16'b0000_0000_0010_0000
  : (A[3:0] == 4'b0110) ? 16'b0000_0000_0100_0000
  : (A[3:0] == 4'b0111) ? 16'b0000_0000_1000_0000
  : (A[3:0] == 4'b1000) ? 16'b0000_0001_0000_0000
  : (A[3:0] == 4'b1001) ? 16'b0000_0010_0000_0000
  : (A[3:0] == 4'b1010) ? 16'b0000_0100_0000_0000
  : (A[3:0] == 4'b1011) ? 16'b0000_1000_0000_0000
  : (A[3:0] == 4'b1100) ? 16'b0001_0000_0000_0000
  : (A[3:0] == 4'b1101) ? 16'b0010_0000_0000_0000
  : (A[3:0] == 4'b1110) ? 16'b0100_0000_0000_0000
  : (A[3:0] == 4'b1111) ? 16'b1000_0000_0000_0000
  : 16'b0000_0000_0000_0000;
endmodule
